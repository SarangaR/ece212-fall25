
module decoder(
    input [1:0] in,
    output reg [3:0] out
);
    //Your code here


endmodule