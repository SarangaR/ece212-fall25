`timescale 1ns/100ps
module xor2_tb();
    //Your code here
    initial begin
        $finish;
    end
endmodule